module interrupt_controller(
	input wire [7:0]int_request,
	input wire irqa,
	
	output wire [7:0]int_no
) ;
reg [31:0]queue1 ;
reg [31:0]queue2 ;


endmodule