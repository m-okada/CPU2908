module xorshift(
	input wire mode,
	input wire clk,
	input [31:0]seed,
	output wire[7:0] rnd
);



endmodule
